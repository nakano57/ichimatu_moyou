localparam HPERIOD = 12'd800;
localparam HFRONT = 12'd16;
localparam HWIDTH = 12'd96;
localparam HBACK = 12'd48;

localparam VPERIOD = 12'd525;
localparam VFRONT = 12'd10;
localparam VWIDTH = 12'd2;
localparam VBACK = 12'd33;
